library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

------------------------------- MEMORY MANAGEMENT UNIT ------------------------------

-- Memory management unit to allow allow a dual port 32 bit wide distributed memory IP core
-- to read and write 16 bit data effectively into only the upper memory region (64 - 128). 

-- MEMORY WRITE: Achieved by first reading an entire 32 bit data segment from the write location, 
-- and modifying either the upper or lower 16 bits of read data to the desired data to be written 
-- based upon the LSB of the write address. This is then written to the desired address.

-- MEMORY READ: Read 32 bit value from data at desired read location, and return to the processor
-- either the upper or lower half of this data dependent upon the LSB of the modified read address.
-- Read address is generated by tagging the MSB of the shortened read address with a '1' to ensure
-- only reading/writing the upper half of memory.

-- INSTRUCTION READ: MIA generated by control unit based upon PC is first shortened by removing 
-- 2 MSB's. We then tag the MSB with a 0 so that we can only address from 0 to 63. This modified
-- MIA is then passed to the memory core as the instruction address. As this exists on its own port
-- the corresponding output port from the memory returns the 32 bit instruction directly to the control
-- unit

--------------------------------------------------------------------------------------

entity MMU is
    Port ( ------------ TO/FROM PROCESSOR -----------
			  MIA : in  STD_LOGIC_VECTOR (7 downto 0); 				  -- Memory instruction address
           DMEM_RW_ADDRESS : in  STD_LOGIC_VECTOR (15 downto 0); -- Desired address to read/write to in DMEM
           DMEM_OUT_TOPROC : out  STD_LOGIC_VECTOR (15 downto 0);-- Data out from the memory core to the processing unit
           OEn : in  STD_LOGIC; -- Write enable signal to Output Reg/ memory core
           DMEM_IN_FROMPROC : in  STD_LOGIC_VECTOR (15 downto 0);-- Data to store into the data memory from the processing unit
			  -------------- TO/FROM DMEM --------------
           INST_ADDRESS : out  STD_LOGIC_VECTOR (6 downto 0);    -- Modified MIA address, to retrieve next instruction from lower half of mem
			  DATA_ADDRESS : out STD_LOGIC_VECTOR(6 downto 0);  	  -- Modified DATA address, to retrieve data from upper half of memory
           DMEM_DATA_TOWRITE : out  STD_LOGIC_VECTOR (31 downto 0); -- Modified data to write to processor, using upper/lower half of data at write location
           DMEM_DATA_READOUT : in  STD_LOGIC_VECTOR (31 downto 0); -- Data read in from the memory
           DMEM_WEn : out  STD_LOGIC; 									  -- Actual Write enable signal to Output Reg/ memory core, piped from OEn input port
			  ----------------- TO/FROM MMIO ----------------
           MMIO_DATA : out  STD_LOGIC_VECTOR (15 downto 0);
           MMIO_WEn : out  STD_LOGIC;
			  PB_IN : in STD_LOGIC);
end MMU;

architecture Behavioral of MMU is
	-- Modified MIA address
	signal MIA_Short : STD_LOGIC_VECTOR(6 downto 0);
	-- Modified data read/write address
	signal DMEM_RWA_Short : STD_LOGIC_VECTOR(6 downto 0);
	-- Temporary signal for storing correctly formed data packet for write address
	signal DMEM_IN_internal : STD_LOGIC_VECTOR(31 downto 0);
	-- Bus to store STD_LOGIC signal from pushbutton into, so processor can read expected 16 bit value
	signal PB_IN_bus : STD_LOGIC_VECTOR(15 downto 0);
begin

-- Throw away the 2 most significant bits, down to 6 bits, between 0 and 63
	MIA_Short(5 downto 0)  <= MIA(5 downto 0);

-- We need to tag with a 0 to address lower half of memory (0 - 63)
	MIA_Short(6) <= '0';

-- Set instruction address to the modified MIA bus value
	INST_ADDRESS <= MIA_Short;
	
-------------- READ -------------------

-- Pushbutton connection. Upper 15 bits of this address are set to 0.
-- The LSB is set to the bit from pushbutton, so a pressed button returns h0001.
	PB_IN_bus(15 downto 1) <= (others => '0');
	PB_IN_bus(0) <= PB_IN;

-- Ignore upper bits of desired memory read address as address lines to dual port memory
-- are only 7 bits wide.
	DMEM_RWA_Short(5 downto 0) <= DMEM_RW_ADDRESS(5 downto 0);

-- Tag the memory address for read/write with a 1 to address the upper half of memory always.
	DMEM_RWA_Short(6) <= '1';
	
-- Set 16 bit data output to processor equal to either the upper or lower half of the 32 bit 
-- data at memory read location dependent upon LSB of read address
	DMEM_OUT_TOPROC <=
		PB_IN_bus when DMEM_RW_ADDRESS = "0000000111110000" else
		DMEM_DATA_READOUT(31 downto 16) when DMEM_RWA_Short(0) = '1' else
		DMEM_DATA_READOUT(15 downto 0) when DMEM_RWA_Short(0) = '0' else
		"0000000000000000";
		
-- Set data address line to memory to modified Read/Write address
DATA_ADDRESS <= DMEM_RWA_Short;

------------ WRITE -------------------

-- Pass through Write enable signal generated by FSM to core and to output register.
DMEM_WEn <= OEn;
MMIO_WEn <= OEn;

-- Set upper half of data value to write to upper half of memory location
DMEM_IN_internal(31 downto 16) <= 
		DMEM_DATA_READOUT(31 downto 16) when DMEM_RWA_Short(0) = '0' and OEn = '1' else
		DMEM_IN_FROMPROC;

-- Set lower half of data value to write to lower half of memory location
DMEM_IN_internal(15 downto 0) <= 
		DMEM_DATA_READOUT(15 downto 0) when DMEM_RWA_Short(0) = '1' and OEn = '1' else
		DMEM_IN_FROMPROC;

-- Set data to write to dual port memory to modified write data
DMEM_DATA_TOWRITE <= DMEM_IN_internal;

-- Set value to output to LED register to 16 bit data from processor when write address
MMIO_DATA <=
		DMEM_IN_FROMPROC when DMEM_RW_ADDRESS = "0000000111111000" else
		"0000000000000000";

end Behavioral;

